module clk(
    input clk,
    output new_clk
);

assign new_clk=clk;

endmodule